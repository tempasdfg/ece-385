module is_wall ( input [9:0] Boy_X_Pos, Boy_Y_Pos,
					  output logic is_wall0, is_wall1, is_wall2, is_wall3, is_wall4, is_wall5, is_wall6
					 )
	logic 